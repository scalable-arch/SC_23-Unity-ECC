module GFEXP(a, b);
  input [7:0] a;
  output [7:0] b;

  /*
    GF(2^8)
    primitive polynomial : x^8 + x6 + x^4 + x^3 + x^2 + x + 1 => Unity ECC와 같다.
    a = a^n
    b = n
  */
  
  reg [7:0] binv;
  always_comb
      case (a)
        8'b0000_0000:  binv = 8'd0; // a=a^0 => 0
        8'b0000_0010:  binv = 8'd1; // a=a^1 => 1
        8'b0000_0100:  binv = 8'd2; // a=a^2 => 2
        8'b0000_1000:  binv = 8'd3; 
        8'b0001_0000:  binv = 8'd4; 
        8'b0010_0000:  binv = 8'd5; 
        8'b0100_0000:  binv = 8'd6; 
        8'b1000_0000:  binv = 8'd7; 
        8'b0101_1111:  binv = 8'd8; 
        8'b1011_1110:  binv = 8'd9; 
        8'b0010_0011:  binv = 8'd10;
        8'b0100_0110:  binv = 8'd11;
        8'b1000_1100:  binv = 8'd12;
        8'b0100_0111:  binv = 8'd13;
        8'b1000_1110:  binv = 8'd14;
        8'b0100_0011:  binv = 8'd15;
        8'b1000_0110:  binv = 8'd16;
        8'b0101_0011:  binv = 8'd17;
        8'b1010_0110:  binv = 8'd18;
        8'b0001_0011:  binv = 8'd19;
        8'b0010_0110:  binv = 8'd20;
        8'b0100_1100:  binv = 8'd21;
        8'b1001_1000:  binv = 8'd22;
        8'b0110_1111:  binv = 8'd23;
        8'b1101_1110:  binv = 8'd24;
        8'b1110_0011:  binv = 8'd25;
        8'b1001_1001:  binv = 8'd26;
        8'b0110_1101:  binv = 8'd27;
        8'b1101_1010:  binv = 8'd28;
        8'b1110_1011:  binv = 8'd29;
        8'b1000_1001:  binv = 8'd30;
        8'b0100_1101:  binv = 8'd31;
        8'b1001_1010:  binv = 8'd32;
        8'b0110_1011:  binv = 8'd33;
        8'b1101_0110:  binv = 8'd34;
        8'b1111_0011:  binv = 8'd35;
        8'b1011_1001:  binv = 8'd36;
        8'b0010_1101:  binv = 8'd37;
        8'b0101_1010:  binv = 8'd38;
        8'b1011_0100:  binv = 8'd39;
        8'b0011_0111:  binv = 8'd40;
        8'b0110_1110:  binv = 8'd41;
        8'b1101_1100:  binv = 8'd42;
        8'b1110_0111:  binv = 8'd43;
        8'b1001_0001:  binv = 8'd44;
        8'b0111_1101:  binv = 8'd45;
        8'b1111_1010:  binv = 8'd46;
        8'b1010_1011:  binv = 8'd47;
        8'b0000_1001:  binv = 8'd48;
        8'b0001_0010:  binv = 8'd49;
        8'b0010_0100:  binv = 8'd50;
        8'b0100_1000:  binv = 8'd51;
        8'b1001_0000:  binv = 8'd52;
        8'b0111_1111:  binv = 8'd53;
        8'b1111_1110:  binv = 8'd54;
        8'b1010_0011:  binv = 8'd55;
        8'b0001_1001:  binv = 8'd56;
        8'b0011_0010:  binv = 8'd57;
        8'b0110_0100:  binv = 8'd58;
        8'b1100_1000:  binv = 8'd59;
        8'b1100_1111:  binv = 8'd60;
        8'b1100_0001:  binv = 8'd61;
        8'b1101_1101:  binv = 8'd62;
        8'b1110_0101:  binv = 8'd63;
        8'b1001_0101:  binv = 8'd64;
        8'b0111_0101:  binv = 8'd65;
        8'b1110_1010:  binv = 8'd66;
        8'b1000_1011:  binv = 8'd67;
        8'b0100_1001:  binv = 8'd68;
        8'b1001_0010:  binv = 8'd69;
        8'b0111_1011:  binv = 8'd70;
        8'b1111_0110:  binv = 8'd71;
        8'b1011_0011:  binv = 8'd72;
        8'b0011_1001:  binv = 8'd73;
        8'b0111_0010:  binv = 8'd74;
        8'b1110_0100:  binv = 8'd75;
        8'b1001_0111:  binv = 8'd76;
        8'b0111_0001:  binv = 8'd77;
        8'b1110_0010:  binv = 8'd78;
        8'b1001_1011:  binv = 8'd79;
        8'b0110_1001:  binv = 8'd80;
        8'b1101_0010:  binv = 8'd81;
        8'b1111_1011:  binv = 8'd82;
        8'b1010_1001:  binv = 8'd83;
        8'b0000_1101:  binv = 8'd84;
        8'b0001_1010:  binv = 8'd85;
        8'b0011_0100:  binv = 8'd86;
        8'b0110_1000:  binv = 8'd87;
        8'b1101_0000:  binv = 8'd88;
        8'b1111_1111:  binv = 8'd89;
        8'b1010_0001:  binv = 8'd90;
        8'b0001_1101:  binv = 8'd91;
        8'b0011_1010:  binv = 8'd92;
        8'b0111_0100:  binv = 8'd93;
        8'b1110_1000:  binv = 8'd94;
        8'b1000_1111:  binv = 8'd95;
        8'b0100_0001:  binv = 8'd96;
        8'b1000_0010:  binv = 8'd97;
        8'b0101_1011:  binv = 8'd98;
        8'b1011_0110:  binv = 8'd99;
        8'b0011_0011:  binv = 8'd100;
        8'b0110_0110:  binv = 8'd101;
        8'b1100_1100:  binv = 8'd102;
        8'b1100_0111:  binv = 8'd103;
        8'b1101_0001:  binv = 8'd104;
        8'b1111_1101:  binv = 8'd105;
        8'b1010_0101:  binv = 8'd106;
        8'b0001_0101:  binv = 8'd107;
        8'b0010_1010:  binv = 8'd108;
        8'b0101_0100:  binv = 8'd109;
        8'b1010_1000:  binv = 8'd110;
        8'b0000_1111:  binv = 8'd111;
        8'b0001_1110:  binv = 8'd112;
        8'b0011_1100:  binv = 8'd113;
        8'b0111_1000:  binv = 8'd114;
        8'b1111_0000:  binv = 8'd115;
        8'b1011_1111:  binv = 8'd116;
        8'b0010_0001:  binv = 8'd117;
        8'b0100_0010:  binv = 8'd118;
        8'b1000_0100:  binv = 8'd119;
        8'b0101_0111:  binv = 8'd120;
        8'b1010_1110:  binv = 8'd121;
        8'b0000_0011:  binv = 8'd122;
        8'b0000_0110:  binv = 8'd123;
        8'b0000_1100:  binv = 8'd124;
        8'b0001_1000:  binv = 8'd125;
        8'b0011_0000:  binv = 8'd126;
        8'b0110_0000:  binv = 8'd127;
        8'b1100_0000:  binv = 8'd128;
        8'b1101_1111:  binv = 8'd129;
        8'b1110_0001:  binv = 8'd130;
        8'b1001_1101:  binv = 8'd131;
        8'b0110_0101:  binv = 8'd132;
        8'b1100_1010:  binv = 8'd133;
        8'b1100_1011:  binv = 8'd134;
        8'b1100_1001:  binv = 8'd135;
        8'b1100_1101:  binv = 8'd136;
        8'b1100_0101:  binv = 8'd137;
        8'b1101_0101:  binv = 8'd138;
        8'b1111_0101:  binv = 8'd139;
        8'b1011_0101:  binv = 8'd140;
        8'b0011_0101:  binv = 8'd141;
        8'b0110_1010:  binv = 8'd142;
        8'b1101_0100:  binv = 8'd143;
        8'b1111_0111:  binv = 8'd144;
        8'b1011_0001:  binv = 8'd145;
        8'b0011_1101:  binv = 8'd146;
        8'b0111_1010:  binv = 8'd147;
        8'b1111_0100:  binv = 8'd148;
        8'b1011_0111:  binv = 8'd149;
        8'b0011_0001:  binv = 8'd150;
        8'b0110_0010:  binv = 8'd151;
        8'b1100_0100:  binv = 8'd152;
        8'b1101_0111:  binv = 8'd153;
        8'b1111_0001:  binv = 8'd154;
        8'b1011_1101:  binv = 8'd155;
        8'b0010_0101:  binv = 8'd156;
        8'b0100_1010:  binv = 8'd157;
        8'b1001_0100:  binv = 8'd158;
        8'b0111_0111:  binv = 8'd159;
        8'b1110_1110:  binv = 8'd160;
        8'b1000_0011:  binv = 8'd161;
        8'b0101_1001:  binv = 8'd162;
        8'b1011_0010:  binv = 8'd163;
        8'b0011_1011:  binv = 8'd164;
        8'b0111_0110:  binv = 8'd165;
        8'b1110_1100:  binv = 8'd166;
        8'b1000_0111:  binv = 8'd167;
        8'b0101_0001:  binv = 8'd168;
        8'b1010_0010:  binv = 8'd169;
        8'b0001_1011:  binv = 8'd170;
        8'b0011_0110:  binv = 8'd171;
        8'b0110_1100:  binv = 8'd172;
        8'b1101_1000:  binv = 8'd173;
        8'b1110_1111:  binv = 8'd174;
        8'b1000_0001:  binv = 8'd175;
        8'b0101_1101:  binv = 8'd176;
        8'b1011_1010:  binv = 8'd177;
        8'b0010_1011:  binv = 8'd178;
        8'b0101_0110:  binv = 8'd179;
        8'b1010_1100:  binv = 8'd180;
        8'b0000_0111:  binv = 8'd181;
        8'b0000_1110:  binv = 8'd182;
        8'b0001_1100:  binv = 8'd183;
        8'b0011_1000:  binv = 8'd184;
        8'b0111_0000:  binv = 8'd185;
        8'b1110_0000:  binv = 8'd186;
        8'b1001_1111:  binv = 8'd187;
        8'b0110_0001:  binv = 8'd188;
        8'b1100_0010:  binv = 8'd189;
        8'b1101_1011:  binv = 8'd190;
        8'b1110_1001:  binv = 8'd191;
        8'b1000_1101:  binv = 8'd192;
        8'b0100_0101:  binv = 8'd193;
        8'b1000_1010:  binv = 8'd194;
        8'b0100_1011:  binv = 8'd195;
        8'b1001_0110:  binv = 8'd196;
        8'b0111_0011:  binv = 8'd197;
        8'b1110_0110:  binv = 8'd198;
        8'b1001_0011:  binv = 8'd199;
        8'b0111_1001:  binv = 8'd200;
        8'b1111_0010:  binv = 8'd201;
        8'b1011_1011:  binv = 8'd202;
        8'b0010_1001:  binv = 8'd203;
        8'b0101_0010:  binv = 8'd204;
        8'b1010_0100:  binv = 8'd205;
        8'b0001_0111:  binv = 8'd206;
        8'b0010_1110:  binv = 8'd207;
        8'b0101_1100:  binv = 8'd208;
        8'b1011_1000:  binv = 8'd209;
        8'b0010_1111:  binv = 8'd210;
        8'b0101_1110:  binv = 8'd211;
        8'b1011_1100:  binv = 8'd212;
        8'b0010_0111:  binv = 8'd213;
        8'b0100_1110:  binv = 8'd214;
        8'b1001_1100:  binv = 8'd215;
        8'b0110_0111:  binv = 8'd216;
        8'b1100_1110:  binv = 8'd217;
        8'b1100_0011:  binv = 8'd218;
        8'b1101_1001:  binv = 8'd219;
        8'b1110_1101:  binv = 8'd220;
        8'b1000_0101:  binv = 8'd221;
        8'b0101_0101:  binv = 8'd222;
        8'b1010_1010:  binv = 8'd223;
        8'b0000_1011:  binv = 8'd224;
        8'b0001_0110:  binv = 8'd225;
        8'b0010_1100:  binv = 8'd226;
        8'b0101_1000:  binv = 8'd227;
        8'b1011_0000:  binv = 8'd228;
        8'b0011_1111:  binv = 8'd229;
        8'b0111_1110:  binv = 8'd230;
        8'b1111_1100:  binv = 8'd231;
        8'b1010_0111:  binv = 8'd232;
        8'b0001_0001:  binv = 8'd233;
        8'b0010_0010:  binv = 8'd234;
        8'b0100_0100:  binv = 8'd235;
        8'b1000_1000:  binv = 8'd236;
        8'b0100_1111:  binv = 8'd237;
        8'b1001_1110:  binv = 8'd238;
        8'b0110_0011:  binv = 8'd239;
        8'b1100_0110:  binv = 8'd240;
        8'b1101_0011:  binv = 8'd241;
        8'b1111_1001:  binv = 8'd242;
        8'b1010_1101:  binv = 8'd243;
        8'b0000_0101:  binv = 8'd244;
        8'b0000_1010:  binv = 8'd245;
        8'b0001_0100:  binv = 8'd246;
        8'b0010_1000:  binv = 8'd247;
        8'b0101_0000:  binv = 8'd248;
        8'b1010_0000:  binv = 8'd249;
        8'b0001_1111:  binv = 8'd250;
        8'b0011_1110:  binv = 8'd251;
        8'b0111_1100:  binv = 8'd252;
        8'b1111_1000:  binv = 8'd253;
        8'b1010_1111:  binv = 8'd254;

      endcase
    assign b = binv;

endmodule


